    NoItem 0NoPath 0NoItem 1NoPath 1NoItem 2NoPath 2NoItem 3NoPath 3NoItem 4NoPath 4NoItem 5NoPath 5NoItem 6NoPath 6NoItem 7NoPath 7NoItem 8NoPath 8NoItem 9NoPath 9               pC�2_    ����?                      �@�2_                               �@�2_                               �@�2_                               �@�2_                                              d       
      $@      4@      Y@      @      $@      Y@����              >@      >@      0@                     �r@      @      Y@      4@     �A@   ����?   ����?   �̬Q@                      �?      $@                              �?    �����	���������	�����������������2D:\DSNetwork\DSN_Structure\usr\bin\KBI20090605.xls                                                                         ��@                 ������.\pRaport9.exe����� �� ��.\pOreolSetTime.exe����� ������.\pOreolVolumeReset.exe
����������.\pOreolSetBlock.exe����� ���������.\pOreolRestart.exepOreolVolumeReset3#E:\Oreol\bin\pOreolVolumeReset3.exeNoItem 6NoPath 6NoItem 7NoPath 7NoItem 8NoPath 8NoItem 9NoPath 9                   4D   A  ���2@  (h0� @              pB   A  ���jk@  (h0� @              �D   A  �>G"@  (h0� @              �C   A  �>GB@  (h0� @              �D   A  �>G"@  (h0� @   �   �  